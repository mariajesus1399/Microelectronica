module contador32bits ( gnd, vdd, enable, clk, reset, mode, D, load, rco, Q);

input gnd, vdd;
input enable;
input clk;
input reset;
output load;
output rco;
input [1:0] mode;
input [3:0] D;
output [31:0] Q;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(mode[1]), .Y(mode_1_bF_buf3) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(mode[1]), .Y(mode_1_bF_buf2) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(mode[1]), .Y(mode_1_bF_buf1) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(mode[1]), .Y(mode_1_bF_buf0) );
	BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(mode[0]), .Y(mode_0_bF_buf3) );
	BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(mode[0]), .Y(mode_0_bF_buf2) );
	BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(mode[0]), .Y(mode_0_bF_buf1) );
	BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(mode[0]), .Y(mode_0_bF_buf0) );
	BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf3) );
	BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf2) );
	BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf1) );
	BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf0) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_373__0_), .Q(\_genblock_contador32bits_v_36_20_0__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_373__1_), .Q(\_genblock_contador32bits_v_36_20_0__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_373__2_), .Q(\_genblock_contador32bits_v_36_20_0__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_373__3_), .Q(\_genblock_contador32bits_v_36_20_0__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_374_), .Q(_0_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .Y(_427_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf3), .Y(_428_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .Y(_429_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_428_), .C(_429_), .Y(_430_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_430_), .Y(_431_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(enable), .Y(_432_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_enable), .B(_432_), .Y(_433_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(op_Q_0_), .Y(_434_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(_434_), .Y(_435_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(op_Q_3_), .Y(_436_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_2_), .Y(_437_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_436_), .Y(_438_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_438_), .C(_433_), .Y(_439_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_439_), .Y(_440_) );
	NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_0_), .C(op_Q_2_), .Y(_441_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_0_), .C(op_Q_2_), .Y(_442_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_442_), .Y(_443_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .Y(_444_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(op_Q_3_), .B(_441_), .Y(_445_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_0_), .Y(_446_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(op_Q_2_), .B(_446_), .C(_436_), .Y(_447_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_447_), .Y(_448_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .Y(_449_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(op_Q_0_), .B(_449_), .Y(_450_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf2), .B(_427_), .C(_429_), .Y(_451_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_451_), .Y(_452_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_452_), .C(_448_), .Y(_453_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .B(_428_), .C(_429_), .Y(_454_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_454_), .Y(_455_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(op_Q_3_), .Y(_456_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_444_), .C(_456_), .Y(_457_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_457_), .C(_453_), .Y(_426_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .B(mode_0_bF_buf1), .Y(_458_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_432_), .Y(_459_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(_458_), .C(_459_), .D(_430_), .Y(_425_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_451_), .Y(_460_) );
	INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_454_), .Y(_461_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_461_), .C(_434_), .Y(_462_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_435_), .Y(_463_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(_434_), .Y(_464_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_463_), .C(_431_), .Y(_465_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .B(_458_), .Y(_466_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_466_), .Y(_467_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_467_), .C(_462_), .Y(_424__0_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_0_), .Y(_468_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(enable), .C(_430_), .Y(_469_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(op_Q_1_), .C(_469_), .Y(_470_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_461_), .C(_468_), .Y(_471_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_466_), .Y(_472_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_472_), .C(_470_), .Y(_424__1_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(enable), .B(op_Q_0_), .Y(_473_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(op_Q_2_), .Y(_474_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_473_), .C(_474_), .Y(_475_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_437_), .B(_473_), .C(_475_), .Y(_476_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_430_), .Y(_477_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_443_), .C(_460_), .Y(_478_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_466_), .C(_461_), .D(_444_), .Y(_479_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_479_), .C(_477_), .Y(_424__2_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_445_), .C(_447_), .Y(_480_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .B(op_Q_0_), .C(op_Q_2_), .Y(_481_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(op_Q_3_), .Y(_482_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_436_), .C(_430_), .Y(_483_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_482_), .C(_483_), .Y(_484_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_466_), .C(_461_), .D(_456_), .Y(_485_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_484_), .C(_485_), .Y(_424__3_) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_424__0_), .Q(op_Q_0_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_424__1_), .Q(op_Q_1_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_424__2_), .Q(op_Q_2_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_424__3_), .Q(op_Q_3_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_425_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_426_), .Q(_genblock_contador32bits_v_36_14_24__op_enable) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(op_Q_0_), .Y(Q[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(op_Q_1_), .Y(Q[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(op_Q_2_), .Y(Q[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(op_Q_3_), .Y(Q[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(Q[4]) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_Q_1_), .Y(Q[5]) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(Q[6]) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(Q[7]) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(Q[8]) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_15_20__op_Q_1_), .Y(Q[9]) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(Q[10]) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(Q[11]) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(Q[12]) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_16_16__op_Q_1_), .Y(Q[13]) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(Q[14]) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(Q[15]) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(Q[16]) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_17_12__op_Q_1_), .Y(Q[17]) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(Q[18]) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(Q[19]) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(Q[20]) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_18_8__op_Q_1_), .Y(Q[21]) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(Q[22]) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(Q[23]) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(Q[24]) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_19_4__op_Q_1_), .Y(Q[25]) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(Q[26]) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(Q[27]) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(Q[28]) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .Y(Q[29]) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(Q[30]) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(Q[31]) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(load) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_undef), .Y(rco) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .Y(_4_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf0), .Y(_5_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .Y(_6_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_4_), .B(_5_), .C(_6_), .Y(_7_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(_8_) );
	INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_enable), .Y(_9_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_14_24__op_rco), .B(_9_), .Y(_10_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_11_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_11_), .Y(_12_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_13_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_14_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_13_), .Y(_15_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_15_), .C(_10_), .Y(_16_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_16_), .Y(_17_) );
	NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_18_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_19_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(_20_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_20_), .Y(_21_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_3_), .B(_18_), .Y(_22_) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_23_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_2_), .B(_23_), .C(_13_), .Y(_24_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_24_), .Y(_25_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .Y(_26_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_0_), .B(_26_), .Y(_27_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf3), .B(_4_), .C(_6_), .Y(_28_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_28_), .Y(_29_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_29_), .C(_25_), .Y(_30_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .B(_5_), .C(_6_), .Y(_31_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_31_), .Y(_32_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_33_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_21_), .C(_33_), .Y(_34_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_34_), .C(_30_), .Y(_3_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .B(mode_0_bF_buf2), .Y(_35_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_9_), .Y(_36_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(_35_), .C(_36_), .D(_7_), .Y(_2_) );
	INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(_37_) );
	INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(_38_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_38_), .C(_11_), .Y(_39_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(_40_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_11_), .Y(_41_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_40_), .C(_8_), .Y(_42_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(_35_), .Y(_43_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_43_), .Y(_44_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .C(_39_), .Y(_1__0_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_45_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_genblock_contador32bits_v_36_14_24__op_enable), .C(_7_), .Y(_46_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_genblock_contador32bits_v_36_14_24__op_Q_1_), .C(_46_), .Y(_47_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_38_), .C(_45_), .Y(_48_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_43_), .Y(_49_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_49_), .C(_47_), .Y(_1__1_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_50_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_51_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_50_), .C(_51_), .Y(_52_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_50_), .C(_52_), .Y(_53_) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_7_), .Y(_54_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_20_), .C(_37_), .Y(_55_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_43_), .C(_38_), .D(_21_), .Y(_56_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_56_), .C(_54_), .Y(_1__2_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_22_), .C(_24_), .Y(_57_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_58_) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_59_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_13_), .C(_7_), .Y(_60_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_59_), .C(_60_), .Y(_61_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_43_), .C(_38_), .D(_33_), .Y(_62_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_61_), .C(_62_), .Y(_1__3_) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_1__0_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_1__1_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_1__2_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1__3_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3_), .Q(_genblock_contador32bits_v_36_14_24__op_rco) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .Y(_66_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf1), .Y(_67_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .Y(_68_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_67_), .C(_68_), .Y(_69_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
	INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_rco), .Y(_71_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_15_20__op_rco), .B(_71_), .Y(_72_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_73_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_73_), .Y(_74_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_75_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_76_) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_75_), .Y(_77_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_77_), .C(_72_), .Y(_78_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_70_), .B(_78_), .Y(_79_) );
	NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_80_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_81_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_81_), .Y(_82_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_82_), .Y(_83_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_3_), .B(_80_), .Y(_84_) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_85_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_2_), .B(_85_), .C(_75_), .Y(_86_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_86_), .Y(_87_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .Y(_88_) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_0_), .B(_88_), .Y(_89_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf0), .B(_66_), .C(_68_), .Y(_90_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .Y(_91_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_91_), .C(_87_), .Y(_92_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .B(_67_), .C(_68_), .Y(_93_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_93_), .Y(_94_) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_95_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_83_), .C(_95_), .Y(_96_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_96_), .C(_92_), .Y(_65_) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .B(mode_0_bF_buf3), .Y(_97_) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_71_), .Y(_98_) );
	OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_97_), .C(_98_), .D(_69_), .Y(_64_) );
	INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_90_), .Y(_99_) );
	INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_100_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .C(_73_), .Y(_101_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_74_), .Y(_102_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_73_), .Y(_103_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_102_), .C(_70_), .Y(_104_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(_97_), .Y(_105_) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_105_), .Y(_106_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_106_), .C(_101_), .Y(_63__0_) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_107_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_genblock_contador32bits_v_36_14_24__op_rco), .C(_69_), .Y(_108_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_genblock_contador32bits_v_36_15_20__op_Q_1_), .C(_108_), .Y(_109_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .C(_107_), .Y(_110_) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_105_), .Y(_111_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_109_), .Y(_63__1_) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_112_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_113_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_112_), .C(_113_), .Y(_114_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_112_), .C(_114_), .Y(_115_) );
	OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_69_), .Y(_116_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_82_), .C(_99_), .Y(_117_) );
	AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_105_), .C(_100_), .D(_83_), .Y(_118_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_118_), .C(_116_), .Y(_63__2_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_84_), .C(_86_), .Y(_119_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_120_) );
	XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_121_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_75_), .C(_69_), .Y(_122_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_121_), .C(_122_), .Y(_123_) );
	AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_105_), .C(_100_), .D(_95_), .Y(_124_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_123_), .C(_124_), .Y(_63__3_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_63__0_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_63__1_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_63__2_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_63__3_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_64_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_65_), .Q(_genblock_contador32bits_v_36_15_20__op_rco) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .Y(_128_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf2), .Y(_129_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .Y(_130_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_129_), .C(_130_), .Y(_131_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_131_), .Y(_132_) );
	INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_rco), .Y(_133_) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_16_16__op_rco), .B(_133_), .Y(_134_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_135_) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_135_), .Y(_136_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_137_) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_138_) );
	OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_137_), .Y(_139_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_136_), .B(_139_), .C(_134_), .Y(_140_) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_140_), .Y(_141_) );
	NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_142_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_143_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_143_), .Y(_144_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_144_), .Y(_145_) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_3_), .B(_142_), .Y(_146_) );
	OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_147_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_2_), .B(_147_), .C(_137_), .Y(_148_) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_148_), .Y(_149_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .Y(_150_) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_0_), .B(_150_), .Y(_151_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf1), .B(_128_), .C(_130_), .Y(_152_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_152_), .Y(_153_) );
	NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_153_), .C(_149_), .Y(_154_) );
	NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .B(_129_), .C(_130_), .Y(_155_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_155_), .Y(_156_) );
	XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_157_) );
	NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_145_), .C(_157_), .Y(_158_) );
	NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_158_), .C(_154_), .Y(_127_) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .B(mode_0_bF_buf0), .Y(_159_) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_133_), .Y(_160_) );
	OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .B(_159_), .C(_160_), .D(_131_), .Y(_126_) );
	INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(_152_), .Y(_161_) );
	INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(_155_), .Y(_162_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_135_), .Y(_163_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(_164_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_135_), .Y(_165_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_164_), .C(_132_), .Y(_166_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_159_), .Y(_167_) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_167_), .Y(_168_) );
	NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_168_), .C(_163_), .Y(_125__0_) );
	XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_169_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_genblock_contador32bits_v_36_15_20__op_rco), .C(_131_), .Y(_170_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_genblock_contador32bits_v_36_16_16__op_Q_1_), .C(_170_), .Y(_171_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_169_), .Y(_172_) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_167_), .Y(_173_) );
	NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_173_), .C(_171_), .Y(_125__1_) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_174_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_175_) );
	OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_174_), .C(_175_), .Y(_176_) );
	OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_174_), .C(_176_), .Y(_177_) );
	OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_131_), .Y(_178_) );
	OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_144_), .C(_161_), .Y(_179_) );
	AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_167_), .C(_162_), .D(_145_), .Y(_180_) );
	NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_180_), .C(_178_), .Y(_125__2_) );
	NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_146_), .C(_148_), .Y(_181_) );
	NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_182_) );
	XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_183_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_137_), .C(_131_), .Y(_184_) );
	OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_183_), .C(_184_), .Y(_185_) );
	AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_167_), .C(_162_), .D(_157_), .Y(_186_) );
	NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_185_), .C(_186_), .Y(_125__3_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_125__0_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_125__1_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_125__2_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_125__3_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_126_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_127_), .Q(_genblock_contador32bits_v_36_16_16__op_rco) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .Y(_190_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf3), .Y(_191_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .Y(_192_) );
	NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_192_), .Y(_193_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
	INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_rco), .Y(_195_) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_17_12__op_rco), .B(_195_), .Y(_196_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_197_) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_197_), .Y(_198_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_199_) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_200_) );
	OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_199_), .Y(_201_) );
	OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_201_), .C(_196_), .Y(_202_) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_202_), .Y(_203_) );
	NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_204_) );
	OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_205_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_205_), .Y(_206_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_206_), .Y(_207_) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_3_), .B(_204_), .Y(_208_) );
	OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_209_) );
	OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_2_), .B(_209_), .C(_199_), .Y(_210_) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_210_), .Y(_211_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .Y(_212_) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_0_), .B(_212_), .Y(_213_) );
	NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf2), .B(_190_), .C(_192_), .Y(_214_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_214_), .Y(_215_) );
	NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_215_), .C(_211_), .Y(_216_) );
	NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .B(_191_), .C(_192_), .Y(_217_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_217_), .Y(_218_) );
	XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_219_) );
	NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_207_), .C(_219_), .Y(_220_) );
	NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_220_), .C(_216_), .Y(_189_) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .B(mode_0_bF_buf1), .Y(_221_) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_195_), .Y(_222_) );
	OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(_221_), .C(_222_), .D(_193_), .Y(_188_) );
	INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(_214_), .Y(_223_) );
	INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_217_), .Y(_224_) );
	OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_224_), .C(_197_), .Y(_225_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_198_), .Y(_226_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_197_), .Y(_227_) );
	OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_226_), .C(_194_), .Y(_228_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .B(_221_), .Y(_229_) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_229_), .Y(_230_) );
	NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_230_), .C(_225_), .Y(_187__0_) );
	XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_231_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_genblock_contador32bits_v_36_16_16__op_rco), .C(_193_), .Y(_232_) );
	OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_genblock_contador32bits_v_36_17_12__op_Q_1_), .C(_232_), .Y(_233_) );
	OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_224_), .C(_231_), .Y(_234_) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_229_), .Y(_235_) );
	NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_235_), .C(_233_), .Y(_187__1_) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_236_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_237_) );
	OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_236_), .C(_237_), .Y(_238_) );
	OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_236_), .C(_238_), .Y(_239_) );
	OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_193_), .Y(_240_) );
	OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_206_), .C(_223_), .Y(_241_) );
	AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_229_), .C(_224_), .D(_207_), .Y(_242_) );
	NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_242_), .C(_240_), .Y(_187__2_) );
	NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_208_), .C(_210_), .Y(_243_) );
	NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_244_) );
	XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_245_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_199_), .C(_193_), .Y(_246_) );
	OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_245_), .C(_246_), .Y(_247_) );
	AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_229_), .C(_224_), .D(_219_), .Y(_248_) );
	NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_247_), .C(_248_), .Y(_187__3_) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_187__0_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_187__1_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_187__2_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_187__3_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_188_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_189_), .Q(_genblock_contador32bits_v_36_17_12__op_rco) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .Y(_252_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf0), .Y(_253_) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .Y(_254_) );
	NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_253_), .C(_254_), .Y(_255_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_255_), .Y(_256_) );
	INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_rco), .Y(_257_) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_18_8__op_rco), .B(_257_), .Y(_258_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_259_) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_259_), .Y(_260_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_261_) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_262_) );
	OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_261_), .Y(_263_) );
	OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_263_), .C(_258_), .Y(_264_) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_256_), .B(_264_), .Y(_265_) );
	NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_266_) );
	OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_267_) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(_267_), .Y(_268_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_268_), .Y(_269_) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_3_), .B(_266_), .Y(_270_) );
	OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_271_) );
	OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_2_), .B(_271_), .C(_261_), .Y(_272_) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_272_), .Y(_273_) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .Y(_274_) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_0_), .B(_274_), .Y(_275_) );
	NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf3), .B(_252_), .C(_254_), .Y(_276_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .Y(_277_) );
	NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_277_), .C(_273_), .Y(_278_) );
	NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .B(_253_), .C(_254_), .Y(_279_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_279_), .Y(_280_) );
	XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_281_) );
	NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_269_), .C(_281_), .Y(_282_) );
	NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_282_), .C(_278_), .Y(_251_) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .B(mode_0_bF_buf2), .Y(_283_) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_257_), .Y(_284_) );
	OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(_283_), .C(_284_), .D(_255_), .Y(_250_) );
	INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(_276_), .Y(_285_) );
	INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(_279_), .Y(_286_) );
	OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_286_), .C(_259_), .Y(_287_) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_260_), .Y(_288_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_259_), .Y(_289_) );
	OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_288_), .C(_256_), .Y(_290_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(_283_), .Y(_291_) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_291_), .Y(_292_) );
	NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_292_), .C(_287_), .Y(_249__0_) );
	XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_293_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_genblock_contador32bits_v_36_17_12__op_rco), .C(_255_), .Y(_294_) );
	OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_genblock_contador32bits_v_36_18_8__op_Q_1_), .C(_294_), .Y(_295_) );
	OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_286_), .C(_293_), .Y(_296_) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_291_), .Y(_297_) );
	NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_297_), .C(_295_), .Y(_249__1_) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_298_) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_299_) );
	OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_298_), .C(_299_), .Y(_300_) );
	OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_298_), .C(_300_), .Y(_301_) );
	OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_255_), .Y(_302_) );
	OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_268_), .C(_285_), .Y(_303_) );
	AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_291_), .C(_286_), .D(_269_), .Y(_304_) );
	NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_304_), .C(_302_), .Y(_249__2_) );
	NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_270_), .C(_272_), .Y(_305_) );
	NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_306_) );
	XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_307_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_261_), .C(_255_), .Y(_308_) );
	OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_257_), .B(_307_), .C(_308_), .Y(_309_) );
	AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_291_), .C(_286_), .D(_281_), .Y(_310_) );
	NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_309_), .C(_310_), .Y(_249__3_) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_249__0_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_249__1_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_249__2_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_249__3_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_250_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_251_), .Q(_genblock_contador32bits_v_36_18_8__op_rco) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .Y(_314_) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf1), .Y(_315_) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .Y(_316_) );
	NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .C(_316_), .Y(_317_) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_317_), .Y(_318_) );
	INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_rco), .Y(_319_) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(\_genblock_contador32bits_v_36_19_4__op_rco), .B(_319_), .Y(_320_) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_321_) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_321_), .Y(_322_) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_323_) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_324_) );
	OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_323_), .Y(_325_) );
	OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_325_), .C(_320_), .Y(_326_) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_318_), .B(_326_), .Y(_327_) );
	NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_328_) );
	OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_329_) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_329_), .Y(_330_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_330_), .Y(_331_) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_3_), .B(_328_), .Y(_332_) );
	OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_333_) );
	OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_2_), .B(_333_), .C(_323_), .Y(_334_) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_334_), .Y(_335_) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .Y(_336_) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_0_), .B(_336_), .Y(_337_) );
	NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf0), .B(_314_), .C(_316_), .Y(_338_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_338_), .Y(_339_) );
	NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_331_), .B(_339_), .C(_335_), .Y(_340_) );
	NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .B(_315_), .C(_316_), .Y(_341_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_341_), .Y(_342_) );
	XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_343_) );
	NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_331_), .C(_343_), .Y(_344_) );
	NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_344_), .C(_340_), .Y(_313_) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf3), .B(mode_0_bF_buf3), .Y(_345_) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_319_), .Y(_346_) );
	OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_345_), .C(_346_), .D(_317_), .Y(_312_) );
	INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_338_), .Y(_347_) );
	INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(_341_), .Y(_348_) );
	OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .C(_321_), .Y(_349_) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_322_), .Y(_350_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_321_), .Y(_351_) );
	OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_350_), .C(_318_), .Y(_352_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(_345_), .Y(_353_) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_353_), .Y(_354_) );
	NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_354_), .C(_349_), .Y(_311__0_) );
	XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_355_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_genblock_contador32bits_v_36_18_8__op_rco), .C(_317_), .Y(_356_) );
	OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_genblock_contador32bits_v_36_19_4__op_Q_1_), .C(_356_), .Y(_357_) );
	OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .C(_355_), .Y(_358_) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_353_), .Y(_359_) );
	NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_359_), .C(_357_), .Y(_311__1_) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_360_) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_361_) );
	OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_360_), .C(_361_), .Y(_362_) );
	OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_360_), .C(_362_), .Y(_363_) );
	OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_317_), .Y(_364_) );
	OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_330_), .C(_347_), .Y(_365_) );
	AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_353_), .C(_348_), .D(_331_), .Y(_366_) );
	NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(_364_), .Y(_311__2_) );
	NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_332_), .C(_334_), .Y(_367_) );
	NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_368_) );
	XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_369_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_323_), .C(_317_), .Y(_370_) );
	OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_369_), .C(_370_), .Y(_371_) );
	AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_353_), .C(_348_), .D(_343_), .Y(_372_) );
	NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .C(_372_), .Y(_311__3_) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_311__0_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_311__1_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_311__2_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_311__3_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_312_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_313_), .Q(_genblock_contador32bits_v_36_19_4__op_rco) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf2), .Y(_375_) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf2), .Y(_376_) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .Y(_377_) );
	NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_376_), .C(_377_), .Y(_378_) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(_378_), .Y(_379_) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_rco), .Y(_380_) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_381_) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_381_), .Y(_382_) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(_383_) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_384_) );
	NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_385_) );
	OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_386_) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_386_), .Y(_387_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_387_), .Y(_388_) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_3_), .B(_385_), .Y(_389_) );
	OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_390_) );
	OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_2_), .B(_390_), .C(_383_), .Y(_391_) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .Y(_392_) );
	NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(mode_0_bF_buf1), .B(_375_), .C(_377_), .Y(_393_) );
	NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf1), .B(_376_), .C(_377_), .Y(_394_) );
	XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(_395_) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(mode_1_bF_buf0), .B(mode_0_bF_buf0), .Y(_396_) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_0_), .B(_380_), .Y(_397_) );
	OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .B(_396_), .C(_397_), .D(_378_), .Y(_374_) );
	INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(_393_), .Y(_398_) );
	INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_394_), .Y(_399_) );
	OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_399_), .C(_381_), .Y(_400_) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_382_), .Y(_401_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_381_), .Y(_402_) );
	OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_401_), .C(_379_), .Y(_403_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_396_), .Y(_404_) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(D[0]), .B(_404_), .Y(_405_) );
	NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_405_), .C(_400_), .Y(_373__0_) );
	XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_406_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_406_), .B(_genblock_contador32bits_v_36_19_4__op_rco), .C(_378_), .Y(_407_) );
	OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_genblock_contador32bits_v_36_20_0__op_Q_1_), .C(_407_), .Y(_408_) );
	OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_399_), .C(_406_), .Y(_409_) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(D[1]), .B(_404_), .Y(_410_) );
	NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(_408_), .Y(_373__1_) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_411_) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_412_) );
	OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_392_), .B(_411_), .C(_412_), .Y(_413_) );
	OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_411_), .C(_413_), .Y(_414_) );
	OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_378_), .Y(_415_) );
	OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_387_), .C(_398_), .Y(_416_) );
	AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(D[2]), .B(_404_), .C(_399_), .D(_388_), .Y(_417_) );
	NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(_415_), .Y(_373__2_) );
	NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_389_), .C(_391_), .Y(_418_) );
	NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_419_) );
	XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(_420_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_383_), .C(_378_), .Y(_421_) );
	OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_420_), .C(_421_), .Y(_422_) );
	AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(D[3]), .B(_404_), .C(_399_), .D(_395_), .Y(_423_) );
	NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_422_), .C(_423_), .Y(_373__3_) );
endmodule
