*** SPICE deck for cell nor3entradas{lay} from library nand3
*** Created on mar. dic. 08, 2020 19:08:54
*** Last revised on mar. dic. 08, 2020 19:34:05
*** Written on mar. dic. 08, 2020 19:34:29 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: nor3entradas{lay}
Mnmos@3 Y A gnd gnd N L=0.4U W=1U AS=6.02P AD=3.353P PS=12.067U PD=10.067U
Mnmos@5 gnd B Y gnd N L=0.4U W=1U AS=3.353P AD=6.02P PS=10.067U PD=12.067U
Mnmos@6 Y C gnd gnd N L=0.4U W=1U AS=6.02P AD=3.353P PS=12.067U PD=10.067U
Mpmos@3 net@54 B net@51 vdd P L=0.4U W=2U AS=5.56P AD=9.56P PS=13.2U PD=21.2U
Mpmos@4 net@51 A vdd vdd P L=0.4U W=2U AS=15.16P AD=5.56P PS=26U PD=13.2U
Mpmos@5 pmos@5_diff-bottom C pmos@5_diff-top vdd P L=0.4U W=2U AS=1.2P AD=1.2P PS=5.2U PD=5.2U

* Spice Code nodes in cell cell 'nor3entradas{lay}'
vdd VDD 0 DC 5    
vinA A 0 pulse (0 5 10n .5n .5n 20n)   
vinB B 0 pulse (0 5 10n .5n .5n 20n) 
vinC C 0 pulse (0 5 10n .5n .5n 20n) 
.MODEL N NMOS  
.MODEL P PMOS    
.TRAN 0 80N   .end 
vdd VDD 0 DC 5     
vinA A 0 pulse (0 5 10n .5n .5n 20n)    
vinB B 0 pulse (0 5 10n .5n .5n 20n)  
vinC C 0 pulse (0 5 10n .5n .5n 20n)  
.MODEL N NMOS   
.MODEL P PMOS     
.TRAN 0 80N   
.end 
vdd VDD 0 DC 5    
vinA A 0 pulse (0 5 10n .5n .5n 20n)   
vinB B 0 pulse (0 5 10n .5n .5n 20n) 
vinC C 0 pulse (0 5 10n .5n .5n 20n) 
.MODEL N NMOS  
.MODEL P PMOS    
.TRAN 0 80N   .end 
.END
