*** SPICE deck for cell nand3{lay} from library compuertas
*** Created on lun. dic. 07, 2020 23:31:33
*** Last revised on mar. dic. 08, 2020 19:32:27
*** Written on mar. dic. 08, 2020 19:35:44 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: nand3{lay}
Mnmos@5 net@95 A gnd gnd N L=0.4U W=1U AS=32.82P AD=5.52P PS=30.2U PD=13.4U
Mnmos@6 net@97 B net@95 gnd N L=0.4U W=1U AS=5.52P AD=5.72P PS=13.4U PD=13.8U
Mnmos@7 Y C net@97 gnd N L=0.4U W=1U AS=5.72P AD=4.095P PS=13.8U PD=9.35U
Mpmos@4 Y A vdd vdd P L=0.4U W=2U AS=6.733P AD=4.095P PS=13.733U PD=9.35U
Mpmos@5 vdd B Y vdd P L=0.4U W=2U AS=4.095P AD=6.733P PS=9.35U PD=13.733U
Mpmos@6 Y C vdd vdd P L=0.4U W=2U AS=6.733P AD=4.095P PS=13.733U PD=9.35U

* Spice Code nodes in cell cell 'nand3{lay}'
vdd VDD 0 DC 5    
vinA A 0 pulse (0 5 10n .5n .5n 20n)   
vinB B 0 pulse (0 5 10n .5n .5n 20n) 
vinC C 0 pulse (0 5 10n .5n .5n 20n) 
.MODEL N NMOS  
.MODEL P PMOS    
.TRAN 0 80N   .end 
.TRAN 0 80N  
.end 
.END
