module contador32bits (enable, clk, reset, mode, D, load, rco, Q);

input enable;
input clk;
input reset;
output load;
output rco;
input [1:0] mode;
input [3:0] D;
output [31:0] Q;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX4 BUFX4_1 ( .A(clk), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_2 ( .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_3 ( .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_4 ( .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_5 ( .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_6 ( .A(clk), .Y(clk_bF_buf0) );
	BUFX2 BUFX2_1 ( .A(mode[1]), .Y(mode_1_bF_buf3) );
	BUFX2 BUFX2_2 ( .A(mode[1]), .Y(mode_1_bF_buf2) );
	BUFX2 BUFX2_3 ( .A(mode[1]), .Y(mode_1_bF_buf1) );
	BUFX2 BUFX2_4 ( .A(mode[1]), .Y(mode_1_bF_buf0) );
	BUFX2 BUFX2_5 ( .A(mode[0]), .Y(mode_0_bF_buf3) );
	BUFX2 BUFX2_6 ( .A(mode[0]), .Y(mode_0_bF_buf2) );
	BUFX2 BUFX2_7 ( .A(mode[0]), .Y(mode_0_bF_buf1) );
	BUFX2 BUFX2_8 ( .A(mode[0]), .Y(mode_0_bF_buf0) );
	BUFX2 BUFX2_9 ( .A(reset), .Y(reset_bF_buf3) );
	BUFX2 BUFX2_10 ( .A(reset), .Y(reset_bF_buf2) );
	BUFX2 BUFX2_11 ( .A(reset), .Y(reset_bF_buf1) );
	BUFX2 BUFX2_12 ( .A(reset), .Y(reset_bF_buf0) );
	AOI21X1 AOI21X1_1 ( .A(_417_), .B(_418_), .C(_386_), .Y(_419_) );
	OAI21X1 OAI21X1_1 ( .A(_416_), .B(_419_), .C(_385_), .Y(_420_) );
	NAND2X1 NAND2X1_1 ( .A(_404_), .B(_393_), .Y(_421_) );
	NAND2X1 NAND2X1_2 ( .A(_392_), .B(_391_), .Y(_422_) );
	AOI22X1 AOI22X1_1 ( .A(D[2]), .B(_409_), .C(_422_), .D(_403_), .Y(_423_) );
	NAND3X1 NAND3X1_1 ( .A(_421_), .B(_423_), .C(_420_), .Y(_379__2_) );
	NAND3X1 NAND3X1_2 ( .A(_395_), .B(_403_), .C(_397_), .Y(_424_) );
	NAND3X1 NAND3X1_3 ( .A(\_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(\_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(\_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_425_) );
	XNOR2X1 XNOR2X1_1 ( .A(_425_), .B(\_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(_426_) );
	AOI21X1 AOI21X1_2 ( .A(_386_), .B(_396_), .C(_384_), .Y(_427_) );
	OAI21X1 OAI21X1_2 ( .A(_386_), .B(_426_), .C(_427_), .Y(_428_) );
	AOI22X1 AOI22X1_2 ( .A(D[3]), .B(_409_), .C(_400_), .D(_404_), .Y(_429_) );
	NAND3X1 NAND3X1_4 ( .A(_424_), .B(_428_), .C(_429_), .Y(_379__3_) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf5), .D(_379__0_), .Q(_genblock_contador32bits_v_36_20_0__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf4), .D(_379__1_), .Q(_genblock_contador32bits_v_36_20_0__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf3), .D(_379__2_), .Q(_genblock_contador32bits_v_36_20_0__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf2), .D(_379__3_), .Q(_genblock_contador32bits_v_36_20_0__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf1), .D(_380_), .Q(_0_) );
	INVX1 INVX1_1 ( .A(mode_1_bF_buf3), .Y(_433_) );
	INVX1 INVX1_2 ( .A(mode_0_bF_buf3), .Y(_434_) );
	INVX1 INVX1_3 ( .A(reset_bF_buf3), .Y(_435_) );
	NAND3X1 NAND3X1_5 ( .A(_433_), .B(_434_), .C(_435_), .Y(_436_) );
	INVX1 INVX1_4 ( .A(_436_), .Y(_437_) );
	INVX1 INVX1_5 ( .A(enable), .Y(_438_) );
	NAND2X1 NAND2X1_3 ( .A(\_genblock_contador32bits_v_36_14_24__op_enable), .B(_438_), .Y(_439_) );
	INVX1 INVX1_6 ( .A(op_Q_0_), .Y(_440_) );
	NAND2X1 NAND2X1_4 ( .A(enable), .B(_440_), .Y(_441_) );
	NAND3X1 NAND3X1_6 ( .A(op_Q_1_), .B(op_Q_2_), .C(op_Q_3_), .Y(_442_) );
	OAI21X1 OAI21X1_3 ( .A(_442_), .B(_441_), .C(_439_), .Y(_443_) );
	NAND2X1 NAND2X1_5 ( .A(_437_), .B(_443_), .Y(_444_) );
	INVX1 INVX1_7 ( .A(op_Q_1_), .Y(_445_) );
	INVX1 INVX1_8 ( .A(op_Q_2_), .Y(_446_) );
	NAND3X1 NAND3X1_7 ( .A(_445_), .B(_440_), .C(_446_), .Y(_447_) );
	OAI21X1 OAI21X1_4 ( .A(op_Q_1_), .B(op_Q_0_), .C(op_Q_2_), .Y(_448_) );
	AND2X2 AND2X2_1 ( .A(_447_), .B(_448_), .Y(_449_) );
	NOR2X1 NOR2X1_1 ( .A(op_Q_1_), .B(op_Q_0_), .Y(_450_) );
	NAND3X1 NAND3X1_8 ( .A(_446_), .B(op_Q_3_), .C(_450_), .Y(_451_) );
	INVX1 INVX1_9 ( .A(op_Q_3_), .Y(_452_) );
	NAND2X1 NAND2X1_6 ( .A(_452_), .B(_447_), .Y(_453_) );
	NAND2X1 NAND2X1_7 ( .A(_451_), .B(_453_), .Y(_454_) );
	NAND2X1 NAND2X1_8 ( .A(op_Q_0_), .B(_445_), .Y(_455_) );
	NAND3X1 NAND3X1_9 ( .A(mode_0_bF_buf2), .B(_433_), .C(_435_), .Y(_456_) );
	NOR2X1 NOR2X1_2 ( .A(_455_), .B(_456_), .Y(_457_) );
	NAND3X1 NAND3X1_10 ( .A(_449_), .B(_457_), .C(_454_), .Y(_458_) );
	INVX1 INVX1_10 ( .A(_450_), .Y(_459_) );
	NAND3X1 NAND3X1_11 ( .A(mode_1_bF_buf2), .B(_434_), .C(_435_), .Y(_460_) );
	NOR2X1 NOR2X1_3 ( .A(_460_), .B(_459_), .Y(_461_) );
	XOR2X1 XOR2X1_1 ( .A(_448_), .B(_452_), .Y(_462_) );
	NAND3X1 NAND3X1_12 ( .A(_449_), .B(_462_), .C(_461_), .Y(_463_) );
	NAND3X1 NAND3X1_13 ( .A(_444_), .B(_463_), .C(_458_), .Y(_432_) );
	NAND2X1 NAND2X1_9 ( .A(mode_1_bF_buf1), .B(mode_0_bF_buf1), .Y(_464_) );
	NAND2X1 NAND2X1_10 ( .A(_0_), .B(_438_), .Y(_465_) );
	OAI22X1 OAI22X1_1 ( .A(reset_bF_buf2), .B(_464_), .C(_465_), .D(_436_), .Y(_431_) );
	INVX1 INVX1_11 ( .A(_456_), .Y(_466_) );
	INVX1 INVX1_12 ( .A(_460_), .Y(_467_) );
	OAI21X1 OAI21X1_5 ( .A(_466_), .B(_467_), .C(_440_), .Y(_468_) );
	INVX1 INVX1_13 ( .A(_441_), .Y(_469_) );
	NOR2X1 NOR2X1_4 ( .A(enable), .B(_440_), .Y(_470_) );
	OAI21X1 OAI21X1_6 ( .A(_470_), .B(_469_), .C(_437_), .Y(_471_) );
	NOR2X1 NOR2X1_5 ( .A(reset_bF_buf1), .B(_464_), .Y(_472_) );
	NAND2X1 NAND2X1_11 ( .A(D[0]), .B(_472_), .Y(_473_) );
	NAND3X1 NAND3X1_14 ( .A(_471_), .B(_473_), .C(_468_), .Y(_430__0_) );
	XNOR2X1 XNOR2X1_2 ( .A(op_Q_1_), .B(op_Q_0_), .Y(_474_) );
	AOI21X1 AOI21X1_3 ( .A(_474_), .B(enable), .C(_436_), .Y(_475_) );
	OAI21X1 OAI21X1_7 ( .A(enable), .B(op_Q_1_), .C(_475_), .Y(_476_) );
	OAI21X1 OAI21X1_8 ( .A(_466_), .B(_467_), .C(_474_), .Y(_477_) );
	NAND2X1 NAND2X1_12 ( .A(D[1]), .B(_472_), .Y(_478_) );
	NAND3X1 NAND3X1_15 ( .A(_478_), .B(_477_), .C(_476_), .Y(_430__1_) );
	NOR2X1 NOR2X1_6 ( .A(enable), .B(_446_), .Y(_479_) );
	OAI21X1 OAI21X1_9 ( .A(_445_), .B(_440_), .C(op_Q_2_), .Y(_480_) );
	NAND3X1 NAND3X1_16 ( .A(op_Q_1_), .B(op_Q_0_), .C(_446_), .Y(_481_) );
	AOI21X1 AOI21X1_4 ( .A(_480_), .B(_481_), .C(_438_), .Y(_482_) );
	OAI21X1 OAI21X1_10 ( .A(_479_), .B(_482_), .C(_437_), .Y(_483_) );
	NAND2X1 NAND2X1_13 ( .A(_467_), .B(_449_), .Y(_484_) );
	NAND2X1 NAND2X1_14 ( .A(_448_), .B(_447_), .Y(_485_) );
	AOI22X1 AOI22X1_3 ( .A(D[2]), .B(_472_), .C(_485_), .D(_466_), .Y(_486_) );
	NAND3X1 NAND3X1_17 ( .A(_484_), .B(_486_), .C(_483_), .Y(_430__2_) );
	NAND3X1 NAND3X1_18 ( .A(_451_), .B(_466_), .C(_453_), .Y(_487_) );
	NAND3X1 NAND3X1_19 ( .A(op_Q_1_), .B(op_Q_0_), .C(op_Q_2_), .Y(_488_) );
	XNOR2X1 XNOR2X1_3 ( .A(_488_), .B(op_Q_3_), .Y(_489_) );
	AOI21X1 AOI21X1_5 ( .A(_438_), .B(_452_), .C(_436_), .Y(_490_) );
	OAI21X1 OAI21X1_11 ( .A(_438_), .B(_489_), .C(_490_), .Y(_491_) );
	AOI22X1 AOI22X1_4 ( .A(D[3]), .B(_472_), .C(_462_), .D(_467_), .Y(_492_) );
	NAND3X1 NAND3X1_20 ( .A(_487_), .B(_491_), .C(_492_), .Y(_430__3_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf0), .D(_430__0_), .Q(op_Q_0_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf5), .D(_430__1_), .Q(op_Q_1_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf4), .D(_430__2_), .Q(op_Q_2_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf3), .D(_430__3_), .Q(op_Q_3_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf2), .D(_431_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf1), .D(_432_), .Q(_genblock_contador32bits_v_36_14_24__op_enable) );
	BUFX2 BUFX2_13 ( .A(op_Q_0_), .Y(Q[0]) );
	BUFX2 BUFX2_14 ( .A(op_Q_1_), .Y(Q[1]) );
	BUFX2 BUFX2_15 ( .A(op_Q_2_), .Y(Q[2]) );
	BUFX2 BUFX2_16 ( .A(op_Q_3_), .Y(Q[3]) );
	BUFX2 BUFX2_17 ( .A(\_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(Q[4]) );
	BUFX2 BUFX2_18 ( .A(\_genblock_contador32bits_v_36_14_24__op_Q_1_), .Y(Q[5]) );
	BUFX2 BUFX2_19 ( .A(\_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(Q[6]) );
	BUFX2 BUFX2_20 ( .A(\_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(Q[7]) );
	BUFX2 BUFX2_21 ( .A(\_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(Q[8]) );
	BUFX2 BUFX2_22 ( .A(\_genblock_contador32bits_v_36_15_20__op_Q_1_), .Y(Q[9]) );
	BUFX2 BUFX2_23 ( .A(\_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(Q[10]) );
	BUFX2 BUFX2_24 ( .A(\_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(Q[11]) );
	BUFX2 BUFX2_25 ( .A(\_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(Q[12]) );
	BUFX2 BUFX2_26 ( .A(\_genblock_contador32bits_v_36_16_16__op_Q_1_), .Y(Q[13]) );
	BUFX2 BUFX2_27 ( .A(\_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(Q[14]) );
	BUFX2 BUFX2_28 ( .A(\_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(Q[15]) );
	BUFX2 BUFX2_29 ( .A(\_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(Q[16]) );
	BUFX2 BUFX2_30 ( .A(\_genblock_contador32bits_v_36_17_12__op_Q_1_), .Y(Q[17]) );
	BUFX2 BUFX2_31 ( .A(\_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(Q[18]) );
	BUFX2 BUFX2_32 ( .A(\_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(Q[19]) );
	BUFX2 BUFX2_33 ( .A(\_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(Q[20]) );
	BUFX2 BUFX2_34 ( .A(\_genblock_contador32bits_v_36_18_8__op_Q_1_), .Y(Q[21]) );
	BUFX2 BUFX2_35 ( .A(\_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(Q[22]) );
	BUFX2 BUFX2_36 ( .A(\_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(Q[23]) );
	BUFX2 BUFX2_37 ( .A(\_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(Q[24]) );
	BUFX2 BUFX2_38 ( .A(\_genblock_contador32bits_v_36_19_4__op_Q_1_), .Y(Q[25]) );
	BUFX2 BUFX2_39 ( .A(\_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(Q[26]) );
	BUFX2 BUFX2_40 ( .A(\_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(Q[27]) );
	BUFX2 BUFX2_41 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(Q[28]) );
	BUFX2 BUFX2_42 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .Y(Q[29]) );
	BUFX2 BUFX2_43 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(Q[30]) );
	BUFX2 BUFX2_44 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(Q[31]) );
	BUFX2 BUFX2_45 ( .A(_0_), .Y(load) );
	BUFX2 BUFX2_46 ( .A(_undef), .Y(rco) );
	INVX1 INVX1_14 ( .A(mode_1_bF_buf0), .Y(_4_) );
	INVX1 INVX1_15 ( .A(mode_0_bF_buf0), .Y(_5_) );
	INVX1 INVX1_16 ( .A(reset_bF_buf0), .Y(_6_) );
	NAND3X1 NAND3X1_21 ( .A(_4_), .B(_5_), .C(_6_), .Y(_7_) );
	INVX1 INVX1_17 ( .A(_7_), .Y(_8_) );
	INVX1 INVX1_18 ( .A(_genblock_contador32bits_v_36_14_24__op_enable), .Y(_9_) );
	NAND2X1 NAND2X1_15 ( .A(\_genblock_contador32bits_v_36_14_24__op_rco), .B(_9_), .Y(_10_) );
	INVX1 INVX1_19 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_11_) );
	NAND2X1 NAND2X1_16 ( .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_11_), .Y(_12_) );
	NAND3X1 NAND3X1_22 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_2_), .C(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_13_) );
	OAI21X1 OAI21X1_12 ( .A(_13_), .B(_12_), .C(_10_), .Y(_14_) );
	NAND2X1 NAND2X1_17 ( .A(_8_), .B(_14_), .Y(_15_) );
	INVX1 INVX1_20 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .Y(_16_) );
	INVX1 INVX1_21 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_17_) );
	NAND3X1 NAND3X1_23 ( .A(_16_), .B(_11_), .C(_17_), .Y(_18_) );
	OAI21X1 OAI21X1_13 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_19_) );
	AND2X2 AND2X2_2 ( .A(_18_), .B(_19_), .Y(_20_) );
	NOR2X1 NOR2X1_7 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_21_) );
	NAND3X1 NAND3X1_24 ( .A(_17_), .B(_genblock_contador32bits_v_36_14_24__op_Q_3_), .C(_21_), .Y(_22_) );
	INVX1 INVX1_22 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_23_) );
	NAND2X1 NAND2X1_18 ( .A(_23_), .B(_18_), .Y(_24_) );
	NAND2X1 NAND2X1_19 ( .A(_22_), .B(_24_), .Y(_25_) );
	NAND2X1 NAND2X1_20 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_0_), .B(_16_), .Y(_26_) );
	NAND3X1 NAND3X1_25 ( .A(mode_0_bF_buf3), .B(_4_), .C(_6_), .Y(_27_) );
	NOR2X1 NOR2X1_8 ( .A(_26_), .B(_27_), .Y(_28_) );
	NAND3X1 NAND3X1_26 ( .A(_20_), .B(_28_), .C(_25_), .Y(_29_) );
	INVX1 INVX1_23 ( .A(_21_), .Y(_30_) );
	NAND3X1 NAND3X1_27 ( .A(mode_1_bF_buf3), .B(_5_), .C(_6_), .Y(_31_) );
	NOR2X1 NOR2X1_9 ( .A(_31_), .B(_30_), .Y(_32_) );
	XOR2X1 XOR2X1_2 ( .A(_19_), .B(_23_), .Y(_33_) );
	NAND3X1 NAND3X1_28 ( .A(_20_), .B(_33_), .C(_32_), .Y(_34_) );
	NAND3X1 NAND3X1_29 ( .A(_15_), .B(_34_), .C(_29_), .Y(_3_) );
	NAND2X1 NAND2X1_21 ( .A(mode_1_bF_buf2), .B(mode_0_bF_buf2), .Y(_35_) );
	NAND2X1 NAND2X1_22 ( .A(_0_), .B(_9_), .Y(_36_) );
	OAI22X1 OAI22X1_2 ( .A(reset_bF_buf3), .B(_35_), .C(_36_), .D(_7_), .Y(_2_) );
	INVX1 INVX1_24 ( .A(_27_), .Y(_37_) );
	INVX1 INVX1_25 ( .A(_31_), .Y(_38_) );
	OAI21X1 OAI21X1_14 ( .A(_37_), .B(_38_), .C(_11_), .Y(_39_) );
	INVX1 INVX1_26 ( .A(_12_), .Y(_40_) );
	NOR2X1 NOR2X1_10 ( .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_11_), .Y(_41_) );
	OAI21X1 OAI21X1_15 ( .A(_41_), .B(_40_), .C(_8_), .Y(_42_) );
	NOR2X1 NOR2X1_11 ( .A(reset_bF_buf2), .B(_35_), .Y(_43_) );
	NAND2X1 NAND2X1_23 ( .A(D[0]), .B(_43_), .Y(_44_) );
	NAND3X1 NAND3X1_30 ( .A(_42_), .B(_44_), .C(_39_), .Y(_1__0_) );
	XNOR2X1 XNOR2X1_4 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .Y(_45_) );
	AOI21X1 AOI21X1_6 ( .A(_45_), .B(_genblock_contador32bits_v_36_14_24__op_enable), .C(_7_), .Y(_46_) );
	OAI21X1 OAI21X1_16 ( .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_genblock_contador32bits_v_36_14_24__op_Q_1_), .C(_46_), .Y(_47_) );
	OAI21X1 OAI21X1_17 ( .A(_37_), .B(_38_), .C(_45_), .Y(_48_) );
	NAND2X1 NAND2X1_24 ( .A(D[1]), .B(_43_), .Y(_49_) );
	NAND3X1 NAND3X1_31 ( .A(_49_), .B(_48_), .C(_47_), .Y(_1__1_) );
	NOR2X1 NOR2X1_12 ( .A(_genblock_contador32bits_v_36_14_24__op_enable), .B(_17_), .Y(_50_) );
	OAI21X1 OAI21X1_18 ( .A(_16_), .B(_11_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_51_) );
	NAND3X1 NAND3X1_32 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_17_), .Y(_52_) );
	AOI21X1 AOI21X1_7 ( .A(_51_), .B(_52_), .C(_9_), .Y(_53_) );
	OAI21X1 OAI21X1_19 ( .A(_50_), .B(_53_), .C(_8_), .Y(_54_) );
	NAND2X1 NAND2X1_25 ( .A(_38_), .B(_20_), .Y(_55_) );
	NAND2X1 NAND2X1_26 ( .A(_19_), .B(_18_), .Y(_56_) );
	AOI22X1 AOI22X1_5 ( .A(D[2]), .B(_43_), .C(_56_), .D(_37_), .Y(_57_) );
	NAND3X1 NAND3X1_33 ( .A(_55_), .B(_57_), .C(_54_), .Y(_1__2_) );
	NAND3X1 NAND3X1_34 ( .A(_22_), .B(_37_), .C(_24_), .Y(_58_) );
	NAND3X1 NAND3X1_35 ( .A(_genblock_contador32bits_v_36_14_24__op_Q_1_), .B(_genblock_contador32bits_v_36_14_24__op_Q_0_), .C(_genblock_contador32bits_v_36_14_24__op_Q_2_), .Y(_59_) );
	XNOR2X1 XNOR2X1_5 ( .A(_59_), .B(_genblock_contador32bits_v_36_14_24__op_Q_3_), .Y(_60_) );
	AOI21X1 AOI21X1_8 ( .A(_9_), .B(_23_), .C(_7_), .Y(_61_) );
	OAI21X1 OAI21X1_20 ( .A(_9_), .B(_60_), .C(_61_), .Y(_62_) );
	AOI22X1 AOI22X1_6 ( .A(D[3]), .B(_43_), .C(_33_), .D(_38_), .Y(_63_) );
	NAND3X1 NAND3X1_36 ( .A(_58_), .B(_62_), .C(_63_), .Y(_1__3_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf0), .D(_1__0_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf5), .D(_1__1_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf4), .D(_1__2_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf3), .D(_1__3_), .Q(_genblock_contador32bits_v_36_14_24__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf2), .D(_2_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf1), .D(_3_), .Q(_genblock_contador32bits_v_36_14_24__op_rco) );
	INVX1 INVX1_27 ( .A(mode_1_bF_buf1), .Y(_67_) );
	INVX1 INVX1_28 ( .A(mode_0_bF_buf1), .Y(_68_) );
	INVX1 INVX1_29 ( .A(reset_bF_buf1), .Y(_69_) );
	NAND3X1 NAND3X1_37 ( .A(_67_), .B(_68_), .C(_69_), .Y(_70_) );
	INVX1 INVX1_30 ( .A(_70_), .Y(_71_) );
	INVX1 INVX1_31 ( .A(_genblock_contador32bits_v_36_14_24__op_rco), .Y(_72_) );
	NAND2X1 NAND2X1_27 ( .A(\_genblock_contador32bits_v_36_15_20__op_rco), .B(_72_), .Y(_73_) );
	INVX1 INVX1_32 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_74_) );
	NAND2X1 NAND2X1_28 ( .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_74_), .Y(_75_) );
	NAND3X1 NAND3X1_38 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_2_), .C(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_76_) );
	OAI21X1 OAI21X1_21 ( .A(_76_), .B(_75_), .C(_73_), .Y(_77_) );
	NAND2X1 NAND2X1_29 ( .A(_71_), .B(_77_), .Y(_78_) );
	INVX1 INVX1_33 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .Y(_79_) );
	INVX1 INVX1_34 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_80_) );
	NAND3X1 NAND3X1_39 ( .A(_79_), .B(_74_), .C(_80_), .Y(_81_) );
	OAI21X1 OAI21X1_22 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_82_) );
	AND2X2 AND2X2_3 ( .A(_81_), .B(_82_), .Y(_83_) );
	NOR2X1 NOR2X1_13 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_84_) );
	NAND3X1 NAND3X1_40 ( .A(_80_), .B(_genblock_contador32bits_v_36_15_20__op_Q_3_), .C(_84_), .Y(_85_) );
	INVX1 INVX1_35 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_86_) );
	NAND2X1 NAND2X1_30 ( .A(_86_), .B(_81_), .Y(_87_) );
	NAND2X1 NAND2X1_31 ( .A(_85_), .B(_87_), .Y(_88_) );
	NAND2X1 NAND2X1_32 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_0_), .B(_79_), .Y(_89_) );
	NAND3X1 NAND3X1_41 ( .A(mode_0_bF_buf0), .B(_67_), .C(_69_), .Y(_90_) );
	NOR2X1 NOR2X1_14 ( .A(_89_), .B(_90_), .Y(_91_) );
	NAND3X1 NAND3X1_42 ( .A(_83_), .B(_91_), .C(_88_), .Y(_92_) );
	INVX1 INVX1_36 ( .A(_84_), .Y(_93_) );
	NAND3X1 NAND3X1_43 ( .A(mode_1_bF_buf0), .B(_68_), .C(_69_), .Y(_94_) );
	NOR2X1 NOR2X1_15 ( .A(_94_), .B(_93_), .Y(_95_) );
	XOR2X1 XOR2X1_3 ( .A(_82_), .B(_86_), .Y(_96_) );
	NAND3X1 NAND3X1_44 ( .A(_83_), .B(_96_), .C(_95_), .Y(_97_) );
	NAND3X1 NAND3X1_45 ( .A(_78_), .B(_97_), .C(_92_), .Y(_66_) );
	NAND2X1 NAND2X1_33 ( .A(mode_1_bF_buf3), .B(mode_0_bF_buf3), .Y(_98_) );
	NAND2X1 NAND2X1_34 ( .A(_0_), .B(_72_), .Y(_99_) );
	OAI22X1 OAI22X1_3 ( .A(reset_bF_buf0), .B(_98_), .C(_99_), .D(_70_), .Y(_65_) );
	INVX1 INVX1_37 ( .A(_90_), .Y(_100_) );
	INVX1 INVX1_38 ( .A(_94_), .Y(_101_) );
	OAI21X1 OAI21X1_23 ( .A(_100_), .B(_101_), .C(_74_), .Y(_102_) );
	INVX1 INVX1_39 ( .A(_75_), .Y(_103_) );
	NOR2X1 NOR2X1_16 ( .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_74_), .Y(_104_) );
	OAI21X1 OAI21X1_24 ( .A(_104_), .B(_103_), .C(_71_), .Y(_105_) );
	NOR2X1 NOR2X1_17 ( .A(reset_bF_buf3), .B(_98_), .Y(_106_) );
	NAND2X1 NAND2X1_35 ( .A(D[0]), .B(_106_), .Y(_107_) );
	NAND3X1 NAND3X1_46 ( .A(_105_), .B(_107_), .C(_102_), .Y(_64__0_) );
	XNOR2X1 XNOR2X1_6 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .Y(_108_) );
	AOI21X1 AOI21X1_9 ( .A(_108_), .B(_genblock_contador32bits_v_36_14_24__op_rco), .C(_70_), .Y(_109_) );
	OAI21X1 OAI21X1_25 ( .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_genblock_contador32bits_v_36_15_20__op_Q_1_), .C(_109_), .Y(_110_) );
	OAI21X1 OAI21X1_26 ( .A(_100_), .B(_101_), .C(_108_), .Y(_111_) );
	NAND2X1 NAND2X1_36 ( .A(D[1]), .B(_106_), .Y(_112_) );
	NAND3X1 NAND3X1_47 ( .A(_112_), .B(_111_), .C(_110_), .Y(_64__1_) );
	NOR2X1 NOR2X1_18 ( .A(_genblock_contador32bits_v_36_14_24__op_rco), .B(_80_), .Y(_113_) );
	OAI21X1 OAI21X1_27 ( .A(_79_), .B(_74_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_114_) );
	NAND3X1 NAND3X1_48 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_80_), .Y(_115_) );
	AOI21X1 AOI21X1_10 ( .A(_114_), .B(_115_), .C(_72_), .Y(_116_) );
	OAI21X1 OAI21X1_28 ( .A(_113_), .B(_116_), .C(_71_), .Y(_117_) );
	NAND2X1 NAND2X1_37 ( .A(_101_), .B(_83_), .Y(_118_) );
	NAND2X1 NAND2X1_38 ( .A(_82_), .B(_81_), .Y(_119_) );
	AOI22X1 AOI22X1_7 ( .A(D[2]), .B(_106_), .C(_119_), .D(_100_), .Y(_120_) );
	NAND3X1 NAND3X1_49 ( .A(_118_), .B(_120_), .C(_117_), .Y(_64__2_) );
	NAND3X1 NAND3X1_50 ( .A(_85_), .B(_100_), .C(_87_), .Y(_121_) );
	NAND3X1 NAND3X1_51 ( .A(_genblock_contador32bits_v_36_15_20__op_Q_1_), .B(_genblock_contador32bits_v_36_15_20__op_Q_0_), .C(_genblock_contador32bits_v_36_15_20__op_Q_2_), .Y(_122_) );
	XNOR2X1 XNOR2X1_7 ( .A(_122_), .B(_genblock_contador32bits_v_36_15_20__op_Q_3_), .Y(_123_) );
	AOI21X1 AOI21X1_11 ( .A(_72_), .B(_86_), .C(_70_), .Y(_124_) );
	OAI21X1 OAI21X1_29 ( .A(_72_), .B(_123_), .C(_124_), .Y(_125_) );
	AOI22X1 AOI22X1_8 ( .A(D[3]), .B(_106_), .C(_96_), .D(_101_), .Y(_126_) );
	NAND3X1 NAND3X1_52 ( .A(_121_), .B(_125_), .C(_126_), .Y(_64__3_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf0), .D(_64__0_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf5), .D(_64__1_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf4), .D(_64__2_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf3), .D(_64__3_), .Q(_genblock_contador32bits_v_36_15_20__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf2), .D(_65_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf1), .D(_66_), .Q(_genblock_contador32bits_v_36_15_20__op_rco) );
	INVX1 INVX1_40 ( .A(mode_1_bF_buf2), .Y(_130_) );
	INVX1 INVX1_41 ( .A(mode_0_bF_buf2), .Y(_131_) );
	INVX1 INVX1_42 ( .A(reset_bF_buf2), .Y(_132_) );
	NAND3X1 NAND3X1_53 ( .A(_130_), .B(_131_), .C(_132_), .Y(_133_) );
	INVX1 INVX1_43 ( .A(_133_), .Y(_134_) );
	INVX1 INVX1_44 ( .A(_genblock_contador32bits_v_36_15_20__op_rco), .Y(_135_) );
	NAND2X1 NAND2X1_39 ( .A(\_genblock_contador32bits_v_36_16_16__op_rco), .B(_135_), .Y(_136_) );
	INVX1 INVX1_45 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_137_) );
	NAND2X1 NAND2X1_40 ( .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_137_), .Y(_138_) );
	NAND3X1 NAND3X1_54 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_2_), .C(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_139_) );
	OAI21X1 OAI21X1_30 ( .A(_139_), .B(_138_), .C(_136_), .Y(_140_) );
	NAND2X1 NAND2X1_41 ( .A(_134_), .B(_140_), .Y(_141_) );
	INVX1 INVX1_46 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .Y(_142_) );
	INVX1 INVX1_47 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_143_) );
	NAND3X1 NAND3X1_55 ( .A(_142_), .B(_137_), .C(_143_), .Y(_144_) );
	OAI21X1 OAI21X1_31 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_145_) );
	AND2X2 AND2X2_4 ( .A(_144_), .B(_145_), .Y(_146_) );
	NOR2X1 NOR2X1_19 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_147_) );
	NAND3X1 NAND3X1_56 ( .A(_143_), .B(_genblock_contador32bits_v_36_16_16__op_Q_3_), .C(_147_), .Y(_148_) );
	INVX1 INVX1_48 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_149_) );
	NAND2X1 NAND2X1_42 ( .A(_149_), .B(_144_), .Y(_150_) );
	NAND2X1 NAND2X1_43 ( .A(_148_), .B(_150_), .Y(_151_) );
	NAND2X1 NAND2X1_44 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_0_), .B(_142_), .Y(_152_) );
	NAND3X1 NAND3X1_57 ( .A(mode_0_bF_buf1), .B(_130_), .C(_132_), .Y(_153_) );
	NOR2X1 NOR2X1_20 ( .A(_152_), .B(_153_), .Y(_154_) );
	NAND3X1 NAND3X1_58 ( .A(_146_), .B(_154_), .C(_151_), .Y(_155_) );
	INVX1 INVX1_49 ( .A(_147_), .Y(_156_) );
	NAND3X1 NAND3X1_59 ( .A(mode_1_bF_buf1), .B(_131_), .C(_132_), .Y(_157_) );
	NOR2X1 NOR2X1_21 ( .A(_157_), .B(_156_), .Y(_158_) );
	XOR2X1 XOR2X1_4 ( .A(_145_), .B(_149_), .Y(_159_) );
	NAND3X1 NAND3X1_60 ( .A(_146_), .B(_159_), .C(_158_), .Y(_160_) );
	NAND3X1 NAND3X1_61 ( .A(_141_), .B(_160_), .C(_155_), .Y(_129_) );
	NAND2X1 NAND2X1_45 ( .A(mode_1_bF_buf0), .B(mode_0_bF_buf0), .Y(_161_) );
	NAND2X1 NAND2X1_46 ( .A(_0_), .B(_135_), .Y(_162_) );
	OAI22X1 OAI22X1_4 ( .A(reset_bF_buf1), .B(_161_), .C(_162_), .D(_133_), .Y(_128_) );
	INVX1 INVX1_50 ( .A(_153_), .Y(_163_) );
	INVX1 INVX1_51 ( .A(_157_), .Y(_164_) );
	OAI21X1 OAI21X1_32 ( .A(_163_), .B(_164_), .C(_137_), .Y(_165_) );
	INVX1 INVX1_52 ( .A(_138_), .Y(_166_) );
	NOR2X1 NOR2X1_22 ( .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_137_), .Y(_167_) );
	OAI21X1 OAI21X1_33 ( .A(_167_), .B(_166_), .C(_134_), .Y(_168_) );
	NOR2X1 NOR2X1_23 ( .A(reset_bF_buf0), .B(_161_), .Y(_169_) );
	NAND2X1 NAND2X1_47 ( .A(D[0]), .B(_169_), .Y(_170_) );
	NAND3X1 NAND3X1_62 ( .A(_168_), .B(_170_), .C(_165_), .Y(_127__0_) );
	XNOR2X1 XNOR2X1_8 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .Y(_171_) );
	AOI21X1 AOI21X1_12 ( .A(_171_), .B(_genblock_contador32bits_v_36_15_20__op_rco), .C(_133_), .Y(_172_) );
	OAI21X1 OAI21X1_34 ( .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_genblock_contador32bits_v_36_16_16__op_Q_1_), .C(_172_), .Y(_173_) );
	OAI21X1 OAI21X1_35 ( .A(_163_), .B(_164_), .C(_171_), .Y(_174_) );
	NAND2X1 NAND2X1_48 ( .A(D[1]), .B(_169_), .Y(_175_) );
	NAND3X1 NAND3X1_63 ( .A(_175_), .B(_174_), .C(_173_), .Y(_127__1_) );
	NOR2X1 NOR2X1_24 ( .A(_genblock_contador32bits_v_36_15_20__op_rco), .B(_143_), .Y(_176_) );
	OAI21X1 OAI21X1_36 ( .A(_142_), .B(_137_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_177_) );
	NAND3X1 NAND3X1_64 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_143_), .Y(_178_) );
	AOI21X1 AOI21X1_13 ( .A(_177_), .B(_178_), .C(_135_), .Y(_179_) );
	OAI21X1 OAI21X1_37 ( .A(_176_), .B(_179_), .C(_134_), .Y(_180_) );
	NAND2X1 NAND2X1_49 ( .A(_164_), .B(_146_), .Y(_181_) );
	NAND2X1 NAND2X1_50 ( .A(_145_), .B(_144_), .Y(_182_) );
	AOI22X1 AOI22X1_9 ( .A(D[2]), .B(_169_), .C(_182_), .D(_163_), .Y(_183_) );
	NAND3X1 NAND3X1_65 ( .A(_181_), .B(_183_), .C(_180_), .Y(_127__2_) );
	NAND3X1 NAND3X1_66 ( .A(_148_), .B(_163_), .C(_150_), .Y(_184_) );
	NAND3X1 NAND3X1_67 ( .A(_genblock_contador32bits_v_36_16_16__op_Q_1_), .B(_genblock_contador32bits_v_36_16_16__op_Q_0_), .C(_genblock_contador32bits_v_36_16_16__op_Q_2_), .Y(_185_) );
	XNOR2X1 XNOR2X1_9 ( .A(_185_), .B(_genblock_contador32bits_v_36_16_16__op_Q_3_), .Y(_186_) );
	AOI21X1 AOI21X1_14 ( .A(_135_), .B(_149_), .C(_133_), .Y(_187_) );
	OAI21X1 OAI21X1_38 ( .A(_135_), .B(_186_), .C(_187_), .Y(_188_) );
	AOI22X1 AOI22X1_10 ( .A(D[3]), .B(_169_), .C(_159_), .D(_164_), .Y(_189_) );
	NAND3X1 NAND3X1_68 ( .A(_184_), .B(_188_), .C(_189_), .Y(_127__3_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(_127__0_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf5), .D(_127__1_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf4), .D(_127__2_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf3), .D(_127__3_), .Q(_genblock_contador32bits_v_36_16_16__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf2), .D(_128_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf1), .D(_129_), .Q(_genblock_contador32bits_v_36_16_16__op_rco) );
	INVX1 INVX1_53 ( .A(mode_1_bF_buf3), .Y(_193_) );
	INVX1 INVX1_54 ( .A(mode_0_bF_buf3), .Y(_194_) );
	INVX1 INVX1_55 ( .A(reset_bF_buf3), .Y(_195_) );
	NAND3X1 NAND3X1_69 ( .A(_193_), .B(_194_), .C(_195_), .Y(_196_) );
	INVX1 INVX1_56 ( .A(_196_), .Y(_197_) );
	INVX1 INVX1_57 ( .A(_genblock_contador32bits_v_36_16_16__op_rco), .Y(_198_) );
	NAND2X1 NAND2X1_51 ( .A(\_genblock_contador32bits_v_36_17_12__op_rco), .B(_198_), .Y(_199_) );
	INVX1 INVX1_58 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_200_) );
	NAND2X1 NAND2X1_52 ( .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_200_), .Y(_201_) );
	NAND3X1 NAND3X1_70 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_2_), .C(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_202_) );
	OAI21X1 OAI21X1_39 ( .A(_202_), .B(_201_), .C(_199_), .Y(_203_) );
	NAND2X1 NAND2X1_53 ( .A(_197_), .B(_203_), .Y(_204_) );
	INVX1 INVX1_59 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .Y(_205_) );
	INVX1 INVX1_60 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_206_) );
	NAND3X1 NAND3X1_71 ( .A(_205_), .B(_200_), .C(_206_), .Y(_207_) );
	OAI21X1 OAI21X1_40 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_208_) );
	AND2X2 AND2X2_5 ( .A(_207_), .B(_208_), .Y(_209_) );
	NOR2X1 NOR2X1_25 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_210_) );
	NAND3X1 NAND3X1_72 ( .A(_206_), .B(_genblock_contador32bits_v_36_17_12__op_Q_3_), .C(_210_), .Y(_211_) );
	INVX1 INVX1_61 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_212_) );
	NAND2X1 NAND2X1_54 ( .A(_212_), .B(_207_), .Y(_213_) );
	NAND2X1 NAND2X1_55 ( .A(_211_), .B(_213_), .Y(_214_) );
	NAND2X1 NAND2X1_56 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_0_), .B(_205_), .Y(_215_) );
	NAND3X1 NAND3X1_73 ( .A(mode_0_bF_buf2), .B(_193_), .C(_195_), .Y(_216_) );
	NOR2X1 NOR2X1_26 ( .A(_215_), .B(_216_), .Y(_217_) );
	NAND3X1 NAND3X1_74 ( .A(_209_), .B(_217_), .C(_214_), .Y(_218_) );
	INVX1 INVX1_62 ( .A(_210_), .Y(_219_) );
	NAND3X1 NAND3X1_75 ( .A(mode_1_bF_buf2), .B(_194_), .C(_195_), .Y(_220_) );
	NOR2X1 NOR2X1_27 ( .A(_220_), .B(_219_), .Y(_221_) );
	XOR2X1 XOR2X1_5 ( .A(_208_), .B(_212_), .Y(_222_) );
	NAND3X1 NAND3X1_76 ( .A(_209_), .B(_222_), .C(_221_), .Y(_223_) );
	NAND3X1 NAND3X1_77 ( .A(_204_), .B(_223_), .C(_218_), .Y(_192_) );
	NAND2X1 NAND2X1_57 ( .A(mode_1_bF_buf1), .B(mode_0_bF_buf1), .Y(_224_) );
	NAND2X1 NAND2X1_58 ( .A(_0_), .B(_198_), .Y(_225_) );
	OAI22X1 OAI22X1_5 ( .A(reset_bF_buf2), .B(_224_), .C(_225_), .D(_196_), .Y(_191_) );
	INVX1 INVX1_63 ( .A(_216_), .Y(_226_) );
	INVX1 INVX1_64 ( .A(_220_), .Y(_227_) );
	OAI21X1 OAI21X1_41 ( .A(_226_), .B(_227_), .C(_200_), .Y(_228_) );
	INVX1 INVX1_65 ( .A(_201_), .Y(_229_) );
	NOR2X1 NOR2X1_28 ( .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_200_), .Y(_230_) );
	OAI21X1 OAI21X1_42 ( .A(_230_), .B(_229_), .C(_197_), .Y(_231_) );
	NOR2X1 NOR2X1_29 ( .A(reset_bF_buf1), .B(_224_), .Y(_232_) );
	NAND2X1 NAND2X1_59 ( .A(D[0]), .B(_232_), .Y(_233_) );
	NAND3X1 NAND3X1_78 ( .A(_231_), .B(_233_), .C(_228_), .Y(_190__0_) );
	XNOR2X1 XNOR2X1_10 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .Y(_234_) );
	AOI21X1 AOI21X1_15 ( .A(_234_), .B(_genblock_contador32bits_v_36_16_16__op_rco), .C(_196_), .Y(_235_) );
	OAI21X1 OAI21X1_43 ( .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_genblock_contador32bits_v_36_17_12__op_Q_1_), .C(_235_), .Y(_236_) );
	OAI21X1 OAI21X1_44 ( .A(_226_), .B(_227_), .C(_234_), .Y(_237_) );
	NAND2X1 NAND2X1_60 ( .A(D[1]), .B(_232_), .Y(_238_) );
	NAND3X1 NAND3X1_79 ( .A(_238_), .B(_237_), .C(_236_), .Y(_190__1_) );
	NOR2X1 NOR2X1_30 ( .A(_genblock_contador32bits_v_36_16_16__op_rco), .B(_206_), .Y(_239_) );
	OAI21X1 OAI21X1_45 ( .A(_205_), .B(_200_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_240_) );
	NAND3X1 NAND3X1_80 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_206_), .Y(_241_) );
	AOI21X1 AOI21X1_16 ( .A(_240_), .B(_241_), .C(_198_), .Y(_242_) );
	OAI21X1 OAI21X1_46 ( .A(_239_), .B(_242_), .C(_197_), .Y(_243_) );
	NAND2X1 NAND2X1_61 ( .A(_227_), .B(_209_), .Y(_244_) );
	NAND2X1 NAND2X1_62 ( .A(_208_), .B(_207_), .Y(_245_) );
	AOI22X1 AOI22X1_11 ( .A(D[2]), .B(_232_), .C(_245_), .D(_226_), .Y(_246_) );
	NAND3X1 NAND3X1_81 ( .A(_244_), .B(_246_), .C(_243_), .Y(_190__2_) );
	NAND3X1 NAND3X1_82 ( .A(_211_), .B(_226_), .C(_213_), .Y(_247_) );
	NAND3X1 NAND3X1_83 ( .A(_genblock_contador32bits_v_36_17_12__op_Q_1_), .B(_genblock_contador32bits_v_36_17_12__op_Q_0_), .C(_genblock_contador32bits_v_36_17_12__op_Q_2_), .Y(_248_) );
	XNOR2X1 XNOR2X1_11 ( .A(_248_), .B(_genblock_contador32bits_v_36_17_12__op_Q_3_), .Y(_249_) );
	AOI21X1 AOI21X1_17 ( .A(_198_), .B(_212_), .C(_196_), .Y(_250_) );
	OAI21X1 OAI21X1_47 ( .A(_198_), .B(_249_), .C(_250_), .Y(_251_) );
	AOI22X1 AOI22X1_12 ( .A(D[3]), .B(_232_), .C(_222_), .D(_227_), .Y(_252_) );
	NAND3X1 NAND3X1_84 ( .A(_247_), .B(_251_), .C(_252_), .Y(_190__3_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf0), .D(_190__0_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf5), .D(_190__1_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf4), .D(_190__2_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf3), .D(_190__3_), .Q(_genblock_contador32bits_v_36_17_12__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf2), .D(_191_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf1), .D(_192_), .Q(_genblock_contador32bits_v_36_17_12__op_rco) );
	INVX1 INVX1_66 ( .A(mode_1_bF_buf0), .Y(_256_) );
	INVX1 INVX1_67 ( .A(mode_0_bF_buf0), .Y(_257_) );
	INVX1 INVX1_68 ( .A(reset_bF_buf0), .Y(_258_) );
	NAND3X1 NAND3X1_85 ( .A(_256_), .B(_257_), .C(_258_), .Y(_259_) );
	INVX1 INVX1_69 ( .A(_259_), .Y(_260_) );
	INVX1 INVX1_70 ( .A(_genblock_contador32bits_v_36_17_12__op_rco), .Y(_261_) );
	NAND2X1 NAND2X1_63 ( .A(\_genblock_contador32bits_v_36_18_8__op_rco), .B(_261_), .Y(_262_) );
	INVX1 INVX1_71 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_263_) );
	NAND2X1 NAND2X1_64 ( .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_263_), .Y(_264_) );
	NAND3X1 NAND3X1_86 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_2_), .C(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_265_) );
	OAI21X1 OAI21X1_48 ( .A(_265_), .B(_264_), .C(_262_), .Y(_266_) );
	NAND2X1 NAND2X1_65 ( .A(_260_), .B(_266_), .Y(_267_) );
	INVX1 INVX1_72 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .Y(_268_) );
	INVX1 INVX1_73 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_269_) );
	NAND3X1 NAND3X1_87 ( .A(_268_), .B(_263_), .C(_269_), .Y(_270_) );
	OAI21X1 OAI21X1_49 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_271_) );
	AND2X2 AND2X2_6 ( .A(_270_), .B(_271_), .Y(_272_) );
	NOR2X1 NOR2X1_31 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_273_) );
	NAND3X1 NAND3X1_88 ( .A(_269_), .B(_genblock_contador32bits_v_36_18_8__op_Q_3_), .C(_273_), .Y(_274_) );
	INVX1 INVX1_74 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_275_) );
	NAND2X1 NAND2X1_66 ( .A(_275_), .B(_270_), .Y(_276_) );
	NAND2X1 NAND2X1_67 ( .A(_274_), .B(_276_), .Y(_277_) );
	NAND2X1 NAND2X1_68 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_0_), .B(_268_), .Y(_278_) );
	NAND3X1 NAND3X1_89 ( .A(mode_0_bF_buf3), .B(_256_), .C(_258_), .Y(_279_) );
	NOR2X1 NOR2X1_32 ( .A(_278_), .B(_279_), .Y(_280_) );
	NAND3X1 NAND3X1_90 ( .A(_272_), .B(_280_), .C(_277_), .Y(_281_) );
	INVX1 INVX1_75 ( .A(_273_), .Y(_282_) );
	NAND3X1 NAND3X1_91 ( .A(mode_1_bF_buf3), .B(_257_), .C(_258_), .Y(_283_) );
	NOR2X1 NOR2X1_33 ( .A(_283_), .B(_282_), .Y(_284_) );
	XOR2X1 XOR2X1_6 ( .A(_271_), .B(_275_), .Y(_285_) );
	NAND3X1 NAND3X1_92 ( .A(_272_), .B(_285_), .C(_284_), .Y(_286_) );
	NAND3X1 NAND3X1_93 ( .A(_267_), .B(_286_), .C(_281_), .Y(_255_) );
	NAND2X1 NAND2X1_69 ( .A(mode_1_bF_buf2), .B(mode_0_bF_buf2), .Y(_287_) );
	NAND2X1 NAND2X1_70 ( .A(_0_), .B(_261_), .Y(_288_) );
	OAI22X1 OAI22X1_6 ( .A(reset_bF_buf3), .B(_287_), .C(_288_), .D(_259_), .Y(_254_) );
	INVX1 INVX1_76 ( .A(_279_), .Y(_289_) );
	INVX1 INVX1_77 ( .A(_283_), .Y(_290_) );
	OAI21X1 OAI21X1_50 ( .A(_289_), .B(_290_), .C(_263_), .Y(_291_) );
	INVX1 INVX1_78 ( .A(_264_), .Y(_292_) );
	NOR2X1 NOR2X1_34 ( .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_263_), .Y(_293_) );
	OAI21X1 OAI21X1_51 ( .A(_293_), .B(_292_), .C(_260_), .Y(_294_) );
	NOR2X1 NOR2X1_35 ( .A(reset_bF_buf2), .B(_287_), .Y(_295_) );
	NAND2X1 NAND2X1_71 ( .A(D[0]), .B(_295_), .Y(_296_) );
	NAND3X1 NAND3X1_94 ( .A(_294_), .B(_296_), .C(_291_), .Y(_253__0_) );
	XNOR2X1 XNOR2X1_12 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .Y(_297_) );
	AOI21X1 AOI21X1_18 ( .A(_297_), .B(_genblock_contador32bits_v_36_17_12__op_rco), .C(_259_), .Y(_298_) );
	OAI21X1 OAI21X1_52 ( .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_genblock_contador32bits_v_36_18_8__op_Q_1_), .C(_298_), .Y(_299_) );
	OAI21X1 OAI21X1_53 ( .A(_289_), .B(_290_), .C(_297_), .Y(_300_) );
	NAND2X1 NAND2X1_72 ( .A(D[1]), .B(_295_), .Y(_301_) );
	NAND3X1 NAND3X1_95 ( .A(_301_), .B(_300_), .C(_299_), .Y(_253__1_) );
	NOR2X1 NOR2X1_36 ( .A(_genblock_contador32bits_v_36_17_12__op_rco), .B(_269_), .Y(_302_) );
	OAI21X1 OAI21X1_54 ( .A(_268_), .B(_263_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_303_) );
	NAND3X1 NAND3X1_96 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_269_), .Y(_304_) );
	AOI21X1 AOI21X1_19 ( .A(_303_), .B(_304_), .C(_261_), .Y(_305_) );
	OAI21X1 OAI21X1_55 ( .A(_302_), .B(_305_), .C(_260_), .Y(_306_) );
	NAND2X1 NAND2X1_73 ( .A(_290_), .B(_272_), .Y(_307_) );
	NAND2X1 NAND2X1_74 ( .A(_271_), .B(_270_), .Y(_308_) );
	AOI22X1 AOI22X1_13 ( .A(D[2]), .B(_295_), .C(_308_), .D(_289_), .Y(_309_) );
	NAND3X1 NAND3X1_97 ( .A(_307_), .B(_309_), .C(_306_), .Y(_253__2_) );
	NAND3X1 NAND3X1_98 ( .A(_274_), .B(_289_), .C(_276_), .Y(_310_) );
	NAND3X1 NAND3X1_99 ( .A(_genblock_contador32bits_v_36_18_8__op_Q_1_), .B(_genblock_contador32bits_v_36_18_8__op_Q_0_), .C(_genblock_contador32bits_v_36_18_8__op_Q_2_), .Y(_311_) );
	XNOR2X1 XNOR2X1_13 ( .A(_311_), .B(_genblock_contador32bits_v_36_18_8__op_Q_3_), .Y(_312_) );
	AOI21X1 AOI21X1_20 ( .A(_261_), .B(_275_), .C(_259_), .Y(_313_) );
	OAI21X1 OAI21X1_56 ( .A(_261_), .B(_312_), .C(_313_), .Y(_314_) );
	AOI22X1 AOI22X1_14 ( .A(D[3]), .B(_295_), .C(_285_), .D(_290_), .Y(_315_) );
	NAND3X1 NAND3X1_100 ( .A(_310_), .B(_314_), .C(_315_), .Y(_253__3_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf0), .D(_253__0_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf5), .D(_253__1_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf4), .D(_253__2_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf3), .D(_253__3_), .Q(_genblock_contador32bits_v_36_18_8__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf2), .D(_254_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf1), .D(_255_), .Q(_genblock_contador32bits_v_36_18_8__op_rco) );
	INVX1 INVX1_79 ( .A(mode_1_bF_buf1), .Y(_319_) );
	INVX1 INVX1_80 ( .A(mode_0_bF_buf1), .Y(_320_) );
	INVX1 INVX1_81 ( .A(reset_bF_buf1), .Y(_321_) );
	NAND3X1 NAND3X1_101 ( .A(_319_), .B(_320_), .C(_321_), .Y(_322_) );
	INVX1 INVX1_82 ( .A(_322_), .Y(_323_) );
	INVX1 INVX1_83 ( .A(_genblock_contador32bits_v_36_18_8__op_rco), .Y(_324_) );
	NAND2X1 NAND2X1_75 ( .A(\_genblock_contador32bits_v_36_19_4__op_rco), .B(_324_), .Y(_325_) );
	INVX1 INVX1_84 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_326_) );
	NAND2X1 NAND2X1_76 ( .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_326_), .Y(_327_) );
	NAND3X1 NAND3X1_102 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_2_), .C(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_328_) );
	OAI21X1 OAI21X1_57 ( .A(_328_), .B(_327_), .C(_325_), .Y(_329_) );
	NAND2X1 NAND2X1_77 ( .A(_323_), .B(_329_), .Y(_330_) );
	INVX1 INVX1_85 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .Y(_331_) );
	INVX1 INVX1_86 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_332_) );
	NAND3X1 NAND3X1_103 ( .A(_331_), .B(_326_), .C(_332_), .Y(_333_) );
	OAI21X1 OAI21X1_58 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_334_) );
	AND2X2 AND2X2_7 ( .A(_333_), .B(_334_), .Y(_335_) );
	NOR2X1 NOR2X1_37 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_336_) );
	NAND3X1 NAND3X1_104 ( .A(_332_), .B(_genblock_contador32bits_v_36_19_4__op_Q_3_), .C(_336_), .Y(_337_) );
	INVX1 INVX1_87 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_338_) );
	NAND2X1 NAND2X1_78 ( .A(_338_), .B(_333_), .Y(_339_) );
	NAND2X1 NAND2X1_79 ( .A(_337_), .B(_339_), .Y(_340_) );
	NAND2X1 NAND2X1_80 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_0_), .B(_331_), .Y(_341_) );
	NAND3X1 NAND3X1_105 ( .A(mode_0_bF_buf0), .B(_319_), .C(_321_), .Y(_342_) );
	NOR2X1 NOR2X1_38 ( .A(_341_), .B(_342_), .Y(_343_) );
	NAND3X1 NAND3X1_106 ( .A(_335_), .B(_343_), .C(_340_), .Y(_344_) );
	INVX1 INVX1_88 ( .A(_336_), .Y(_345_) );
	NAND3X1 NAND3X1_107 ( .A(mode_1_bF_buf0), .B(_320_), .C(_321_), .Y(_346_) );
	NOR2X1 NOR2X1_39 ( .A(_346_), .B(_345_), .Y(_347_) );
	XOR2X1 XOR2X1_7 ( .A(_334_), .B(_338_), .Y(_348_) );
	NAND3X1 NAND3X1_108 ( .A(_335_), .B(_348_), .C(_347_), .Y(_349_) );
	NAND3X1 NAND3X1_109 ( .A(_330_), .B(_349_), .C(_344_), .Y(_318_) );
	NAND2X1 NAND2X1_81 ( .A(mode_1_bF_buf3), .B(mode_0_bF_buf3), .Y(_350_) );
	NAND2X1 NAND2X1_82 ( .A(_0_), .B(_324_), .Y(_351_) );
	OAI22X1 OAI22X1_7 ( .A(reset_bF_buf0), .B(_350_), .C(_351_), .D(_322_), .Y(_317_) );
	INVX1 INVX1_89 ( .A(_342_), .Y(_352_) );
	INVX1 INVX1_90 ( .A(_346_), .Y(_353_) );
	OAI21X1 OAI21X1_59 ( .A(_352_), .B(_353_), .C(_326_), .Y(_354_) );
	INVX1 INVX1_91 ( .A(_327_), .Y(_355_) );
	NOR2X1 NOR2X1_40 ( .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_326_), .Y(_356_) );
	OAI21X1 OAI21X1_60 ( .A(_356_), .B(_355_), .C(_323_), .Y(_357_) );
	NOR2X1 NOR2X1_41 ( .A(reset_bF_buf3), .B(_350_), .Y(_358_) );
	NAND2X1 NAND2X1_83 ( .A(D[0]), .B(_358_), .Y(_359_) );
	NAND3X1 NAND3X1_110 ( .A(_357_), .B(_359_), .C(_354_), .Y(_316__0_) );
	XNOR2X1 XNOR2X1_14 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .Y(_360_) );
	AOI21X1 AOI21X1_21 ( .A(_360_), .B(_genblock_contador32bits_v_36_18_8__op_rco), .C(_322_), .Y(_361_) );
	OAI21X1 OAI21X1_61 ( .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_genblock_contador32bits_v_36_19_4__op_Q_1_), .C(_361_), .Y(_362_) );
	OAI21X1 OAI21X1_62 ( .A(_352_), .B(_353_), .C(_360_), .Y(_363_) );
	NAND2X1 NAND2X1_84 ( .A(D[1]), .B(_358_), .Y(_364_) );
	NAND3X1 NAND3X1_111 ( .A(_364_), .B(_363_), .C(_362_), .Y(_316__1_) );
	NOR2X1 NOR2X1_42 ( .A(_genblock_contador32bits_v_36_18_8__op_rco), .B(_332_), .Y(_365_) );
	OAI21X1 OAI21X1_63 ( .A(_331_), .B(_326_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_366_) );
	NAND3X1 NAND3X1_112 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_332_), .Y(_367_) );
	AOI21X1 AOI21X1_22 ( .A(_366_), .B(_367_), .C(_324_), .Y(_368_) );
	OAI21X1 OAI21X1_64 ( .A(_365_), .B(_368_), .C(_323_), .Y(_369_) );
	NAND2X1 NAND2X1_85 ( .A(_353_), .B(_335_), .Y(_370_) );
	NAND2X1 NAND2X1_86 ( .A(_334_), .B(_333_), .Y(_371_) );
	AOI22X1 AOI22X1_15 ( .A(D[2]), .B(_358_), .C(_371_), .D(_352_), .Y(_372_) );
	NAND3X1 NAND3X1_113 ( .A(_370_), .B(_372_), .C(_369_), .Y(_316__2_) );
	NAND3X1 NAND3X1_114 ( .A(_337_), .B(_352_), .C(_339_), .Y(_373_) );
	NAND3X1 NAND3X1_115 ( .A(_genblock_contador32bits_v_36_19_4__op_Q_1_), .B(_genblock_contador32bits_v_36_19_4__op_Q_0_), .C(_genblock_contador32bits_v_36_19_4__op_Q_2_), .Y(_374_) );
	XNOR2X1 XNOR2X1_15 ( .A(_374_), .B(_genblock_contador32bits_v_36_19_4__op_Q_3_), .Y(_375_) );
	AOI21X1 AOI21X1_23 ( .A(_324_), .B(_338_), .C(_322_), .Y(_376_) );
	OAI21X1 OAI21X1_65 ( .A(_324_), .B(_375_), .C(_376_), .Y(_377_) );
	AOI22X1 AOI22X1_16 ( .A(D[3]), .B(_358_), .C(_348_), .D(_353_), .Y(_378_) );
	NAND3X1 NAND3X1_116 ( .A(_373_), .B(_377_), .C(_378_), .Y(_316__3_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf0), .D(_316__0_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_0_) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf5), .D(_316__1_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_1_) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf4), .D(_316__2_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_2_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf3), .D(_316__3_), .Q(_genblock_contador32bits_v_36_19_4__op_Q_3_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf2), .D(_317_), .Q(_0_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf1), .D(_318_), .Q(_genblock_contador32bits_v_36_19_4__op_rco) );
	INVX1 INVX1_92 ( .A(mode_1_bF_buf2), .Y(_381_) );
	INVX1 INVX1_93 ( .A(mode_0_bF_buf2), .Y(_382_) );
	INVX1 INVX1_94 ( .A(reset_bF_buf2), .Y(_383_) );
	NAND3X1 NAND3X1_117 ( .A(_381_), .B(_382_), .C(_383_), .Y(_384_) );
	INVX1 INVX1_95 ( .A(_384_), .Y(_385_) );
	INVX1 INVX1_96 ( .A(_genblock_contador32bits_v_36_19_4__op_rco), .Y(_386_) );
	INVX1 INVX1_97 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_387_) );
	NAND2X1 NAND2X1_87 ( .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_387_), .Y(_388_) );
	INVX1 INVX1_98 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .Y(_389_) );
	INVX1 INVX1_99 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_390_) );
	NAND3X1 NAND3X1_118 ( .A(_389_), .B(_387_), .C(_390_), .Y(_391_) );
	OAI21X1 OAI21X1_66 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_392_) );
	AND2X2 AND2X2_8 ( .A(_391_), .B(_392_), .Y(_393_) );
	NOR2X1 NOR2X1_43 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_394_) );
	NAND3X1 NAND3X1_119 ( .A(_390_), .B(_genblock_contador32bits_v_36_20_0__op_Q_3_), .C(_394_), .Y(_395_) );
	INVX1 INVX1_100 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_3_), .Y(_396_) );
	NAND2X1 NAND2X1_88 ( .A(_396_), .B(_391_), .Y(_397_) );
	NAND3X1 NAND3X1_120 ( .A(mode_0_bF_buf1), .B(_381_), .C(_383_), .Y(_398_) );
	NAND3X1 NAND3X1_121 ( .A(mode_1_bF_buf1), .B(_382_), .C(_383_), .Y(_399_) );
	XOR2X1 XOR2X1_8 ( .A(_392_), .B(_396_), .Y(_400_) );
	NAND2X1 NAND2X1_89 ( .A(mode_1_bF_buf0), .B(mode_0_bF_buf0), .Y(_401_) );
	NAND2X1 NAND2X1_90 ( .A(_0_), .B(_386_), .Y(_402_) );
	OAI22X1 OAI22X1_8 ( .A(reset_bF_buf1), .B(_401_), .C(_402_), .D(_384_), .Y(_380_) );
	INVX1 INVX1_101 ( .A(_398_), .Y(_403_) );
	INVX1 INVX1_102 ( .A(_399_), .Y(_404_) );
	OAI21X1 OAI21X1_67 ( .A(_403_), .B(_404_), .C(_387_), .Y(_405_) );
	INVX1 INVX1_103 ( .A(_388_), .Y(_406_) );
	NOR2X1 NOR2X1_44 ( .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_387_), .Y(_407_) );
	OAI21X1 OAI21X1_68 ( .A(_407_), .B(_406_), .C(_385_), .Y(_408_) );
	NOR2X1 NOR2X1_45 ( .A(reset_bF_buf0), .B(_401_), .Y(_409_) );
	NAND2X1 NAND2X1_91 ( .A(D[0]), .B(_409_), .Y(_410_) );
	NAND3X1 NAND3X1_122 ( .A(_408_), .B(_410_), .C(_405_), .Y(_379__0_) );
	XNOR2X1 XNOR2X1_16 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .Y(_411_) );
	AOI21X1 AOI21X1_24 ( .A(_411_), .B(_genblock_contador32bits_v_36_19_4__op_rco), .C(_384_), .Y(_412_) );
	OAI21X1 OAI21X1_69 ( .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_genblock_contador32bits_v_36_20_0__op_Q_1_), .C(_412_), .Y(_413_) );
	OAI21X1 OAI21X1_70 ( .A(_403_), .B(_404_), .C(_411_), .Y(_414_) );
	NAND2X1 NAND2X1_92 ( .A(D[1]), .B(_409_), .Y(_415_) );
	NAND3X1 NAND3X1_123 ( .A(_415_), .B(_414_), .C(_413_), .Y(_379__1_) );
	NOR2X1 NOR2X1_46 ( .A(_genblock_contador32bits_v_36_19_4__op_rco), .B(_390_), .Y(_416_) );
	OAI21X1 OAI21X1_71 ( .A(_389_), .B(_387_), .C(_genblock_contador32bits_v_36_20_0__op_Q_2_), .Y(_417_) );
	NAND3X1 NAND3X1_124 ( .A(_genblock_contador32bits_v_36_20_0__op_Q_1_), .B(_genblock_contador32bits_v_36_20_0__op_Q_0_), .C(_390_), .Y(_418_) );
endmodule
